`define NUM_OF_GATES 3
`define NUM_OF_RO 8
`define GATE_DELAY 2
